module seg_display_output (input logic [3:0] number,
            output [7:0] hex
);

    always @(number) begin
        case (number)
            4'b0000: hex[7:0] = 8'b11000000; // 0
            4'b0001: hex[7:0] = 8'b11111001; // 1
            4'b0010: hex[7:0] = 8'b10100100; // 2
            4'b0011: hex[7:0] = 8'b10110000; // 3
            4'b0100: hex[7:0] = 8'b10011001; // 4
            4'b0101: hex[7:0] = 8'b10010010; // 5
            4'b0110: hex[7:0] = 8'b10000010; // 6
            4'b0111: hex[7:0] = 8'b11111000; // 7
            4'b1000: hex[7:0] = 8'b10000000; // 8
            4'b1001: hex[7:0] = 8'b10010000; // 9
            4'b1010: hex[7:0] = 8'b11111111; // Display nothing
            4'b1011: hex[7:0] = 8'b10111111; // -
            4'b1100: hex[7:0] = 8'b10001100; // P
            4'b1101: hex[7:0] = 8'b00101111; // r.
            4'b1110: hex[7:0] = 8'b00000110; // E.
            4'b1111: hex[7:0] = 8'b10001110; // F
            default: hex[7:0] = 8'b01111111; // .
        endcase 
    end
    
endmodule